`timescale 1ns / 1ps
module core(
    input clk,
    input rst_n
    );
 
endmodule
